// Steven Herbst
// sherbst@stanford.edu

`timescale 1ns/1ps

`include "svreal.sv"
`include "msdsl.sv"

`default_nettype none

module tb(
    input wire logic sw_1,
    input wire logic sw_2,
    input wire logic btn_1,
    input wire logic btn_2,
    output wire logic led_1,
    output wire logic led_2,
    output wire logic rgb_led_1,
    output wire logic rgb_led_2,
    inout wire logic pmod_1,
    inout wire logic pmod_2
);
    // Some dummy signals to verify physical connections
    // logic sw_1, sw_2, led_1, led_2, rgb_led_1, rgb_led_2, btn_1, btn_2, pmod_1, pmod_2, rst_1;

    // input is a fixed value
    `MAKE_CONST_REAL(1.0, v_in);

    // output has range range +/- 1.5
    `MAKE_REAL(v_out, 1.5);

    // filter instantiation
    filter #(
        `PASS_REAL(v_in, v_in),
        `PASS_REAL(v_out, v_out)
    ) filter_i (
        .v_in(v_in),
        .v_out(v_out)
    );

endmodule

`default_nettype wire
